module test()
endmodule
