module test()
always@()
begin
end
endmodule

